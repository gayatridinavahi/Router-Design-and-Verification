`include "router_dut.sv"
`include "router_tb.sv"
